--! This is a wrapper to prevent Vivado from flagging illegal recursive instantiation.
--! It is an exact mirror of the MLD, which *should* work at the top level, but doesn't.
-------------------------------------------------------------------------------------
-- mld_v1_top_alt.vhd
-------------------------------------------------------------------------------------
-- Authors:     Maxwell Phillips
-- Copyright:   Ohio Northern University, 2024.
-- License:     GPL v3
-- Description: Generic, configurable, multi-level decoder.
-- Precision:   Any power of 2 >= 4.
-------------------------------------------------------------------------------------
--
-- Returns 2 to the power of the input.
--
-- ! This decoder is dimensioned as `n : 2^n`. 
-- The primary files are dimensioned `lg(n) : n` for convenient use with 
-- (priority) encoders, but this may not be the best solution for all hardware, 
-- thus the existence of this file.
--
-- Requires VHDL-2008.
--
-------------------------------------------------------------------------------------
-- Generics
-------------------------------------------------------------------------------------
--
-- [G_lg_n]: Input length; base 2 logarithm of output length `n`.
--
-- [G_n]: Output length `n`.
--
-- [G_max_lvls]: Maximum depth of the decoder. Minimum 2. The decoder may not
--  necessarily reach this number of levels, depending on the input size.
--  The smallest decoder is a 2:4 decoder, so if [G_max_lvls] is high enough,
--  and the input size is small enough, the number of levels will be < [G_max_lvls].
--  Has the highest priority of any constraint.
--
-- [G_use_gate_optimized]: Boolean. True if gate-level optimized row-column
--  decoders should be used for the base level of the overarching decoder.
--  Default false. The maximum size for a gate-optimized decoder is 5:32. The
--  gate-level decoders generated by this constraint are two-level and row-column.
--  With higher input precisions, it is more efficient to use multi-level methods.
--  If [G_max_lvls] does not permit a base level decoder to be 5:32 or smaller,
--  a function-based decoder will be generated instead.
--
-- [G_use_cascading]: Boolean. True if cascading should be used instead of
--  composition as a method of constructing the multi-level decoder. Default false.
--  Has no effect if [G_max_lvls] is not greater than 2.
--
-------------------------------------------------------------------------------------
-- Ports
-------------------------------------------------------------------------------------
--
-- [input]: Parallel input of [G_lg_n] bits.
--
-- [output]: Parallel output of [G_n] bits, exactly 2^[input]; alternatively:
--  a vector of zeroes with a single high bit at index corresponding to [input].
--
-------------------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.numeric_std_unsigned.all;
  use IEEE.math_real.all;

--! If TerosHDL flags an error that: 'ml_decoder' is not compiled in library 'work'
--! This can be safely ignored. 
library work;
  use work.ml_decoder;

entity mld_top_alt is
  generic (
    G_n                    : natural := 6;        --! total input width
    G_2_pow_n              : natural := 2 ** G_n; --! total output width
    G_max_lvls             : natural := 2;        --! maximum depth of the encoder
    G_use_gate_optimized   : boolean := true;     --! whether to use gate-level optimized SLDs at the base level
    G_use_cascading        : boolean := false     --! whether to use cascading instead of composition
  );
  port (
    input  : in    std_logic_vector(G_n - 1 downto 0);
    output : out   std_logic_vector(G_2_pow_n - 1 downto 0)
  );
end mld_top_alt;

architecture behavioral of mld_top_alt is

begin

  inst : entity work.ml_decoder(behavioral)
    generic map (
      G_n                    => G_2_pow_n,
      G_lg_n                 => G_n,
      G_max_lvls             => G_max_lvls,
      G_use_gate_optimized   => G_use_gate_optimized,
      G_use_cascading        => G_use_cascading
    )
    port map (
      input  => input,
      output => output
    );

end architecture behavioral;