-------------------------------------------------------------------------------------
-- mld_v1.vhd
-------------------------------------------------------------------------------------
-- Authors:     Maxwell Phillips
-- Copyright:   Ohio Northern University, 2024.
-- License:     GPL v3
-- Description: Generic, configurable, multi-level decoder.
-- Precision:   Any power of 2 >= 4.
-------------------------------------------------------------------------------------
--
-- Returns 2 to the power of the input.
--
-- ! This decoder is dimensioned as `lg(n) : n`, not `n : 2^n`.
-- It is intentionally designed to complement a(n) (priority) encoder.
--
-- Requires VHDL-2008.
--
-------------------------------------------------------------------------------------
-- Generics
-------------------------------------------------------------------------------------
--
-- [G_lg_n]: Input length; base 2 logarithm of output length `n`.
--
-- [G_n]: Output length `n`.
--
-- [G_max_lvls]: Maximum depth of the decoder. Minimum 2. The decoder may not
--  necessarily reach this number of levels, depending on the input size.
--  The smallest decoder is a 2:4 decoder, so if [G_max_lvls] is high enough,
--  and the input size is small enough, the number of levels will be < [G_max_lvls].
--  Has the highest priority of any constraint.
--
-- [G_use_gate_optimized]: Boolean. True if gate-level optimized row-column
--  decoders should be used for the base level of the overarching decoder.
--  Default false. The maximum size for a gate-optimized decoder is 5:32. The
--  gate-level decoders generated by this constraint are two-level and row-column.
--  With higher input precisions, it is more efficient to use multi-level methods.
--  If [G_max_lvls] does not permit a base level decoder to be 5:32 or smaller,
--  a function-based decoder will be generated instead.
--
-- [G_use_cascading]: Boolean. True if cascading should be used instead of
--  composition as a method of constructing the multi-level decoder. Default false.
--  Has no effect if [G_max_lvls] is not greater than 2.
--
-------------------------------------------------------------------------------------
-- Ports
-------------------------------------------------------------------------------------
--
-- [input]: Parallel input of [G_lg_n] bits.
--
-- [output]: Parallel output of [G_n] bits, exactly 2^[input]; alternatively:
--  a vector of zeroes with a single high bit at index corresponding to [input].
--
-------------------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.numeric_std_unsigned.all;
  use IEEE.math_real.all;

entity ml_decoder is
  generic (
    G_n                    : natural := 64;                              --! total output width
    G_lg_n                 : natural := natural(round(log2(real(G_n)))); --! total input width
    G_max_lvls             : natural := 2;                               --! maximum depth of the encoder
    G_use_gate_optimized   : boolean := false;                           --! whether to use gate-level optimized SLDs at the base level
    G_use_cascading        : boolean := false                            --! whether to use cascading instead of composition
  );
  port (
    input  : in    std_logic_vector(G_lg_n - 1 downto 0);
    output : out   std_logic_vector(G_n - 1 downto 0)
  );
end ml_decoder;

architecture behavioral of ml_decoder is

  -- shorthand function to calculate the size of a signal in bits

  function lg (arg: natural) return natural is begin

    return natural(round(log2(real(arg))));

  end function;

  -- * Components

  component ml_decoder is
    generic (
      G_n                    : natural;
      G_lg_n                 : natural;
      G_max_lvls             : natural;
      G_use_gate_optimized   : boolean;
      G_use_cascading        : boolean
    );
    port (
      input  : in    std_logic_vector(G_lg_n - 1 downto 0);
      output : out   std_logic_vector(G_n - 1 downto 0)
    );
  end component;

begin

  -- this implementation works by decrementing [G_max_lvls] each time a level is instantiated.
  -- this block determines if another sub-level should be generated,
  --  or if the base level of single-level decoders should be generated instead.
  determine_level :
  if G_max_lvls > 1 generate -- generate another level

    -- determine whether to use composite or cascading structure.
    -- when [G_max_lvls] is 1, a single-level decoder is generated (this is the base case).
    -- when [G_max_lvls] is 2, composition is used, regardless of the value of [G_use_cascading].
    --  the result would be the same, but it makes more sense to do this.
    -- when [G_max_lvls] is 3 or higher, a composed or cascaded decoder is generated with
    --  a number of levels less than or equal to [G_max_lvls].
    determine_encoder_type :
    if (not G_use_cascading) or (G_max_lvls < 3) generate

      -- "coarse" decoder handles "columns"
      -- "fine" decoder handles "rows"

      -- * Configuration "Variables"
      constant f    : natural := natural(round(2 ** ceil(log2(sqrt(real(G_n))))));  -- fine decoder output width
      constant lg_f : natural := lg(f);                                             -- fine decoder input width
      constant c    : natural := G_n / f;                                           -- coarse decoder output width
      constant lg_c : natural := lg(c);                                             -- coarse decoder input width

      signal c_input  : std_logic_vector(lg_c - 1 downto 0);  -- coarse decoder input
      signal c_output : std_logic_vector(c - 1 downto 0);     -- coarse decoder output
      signal f_input  : std_logic_vector(lg_f - 1 downto 0);  -- fine decoder input
      signal f_output : std_logic_vector(f - 1 downto 0);     -- fine decoder output

    begin

      c_input <= input(G_lg_n - 1 downto lg_f);
      f_input <= input(lg_f - 1 downto 0);

      coarse_encoder : ml_decoder
        generic map (
          G_n                    => c,
          G_lg_n                 => lg_c,
          G_max_lvls             => (G_max_lvls - 1),
          G_use_gate_optimized   => G_use_gate_optimized,
          G_use_cascading        => G_use_cascading
        )
        port map (
          input  => c_input,
          output => c_output
        );

      fine_encoder : ml_decoder
        generic map (
          G_n                    => f,
          G_lg_n                 => lg_f,
          G_max_lvls             => (G_max_lvls - 1),
          G_use_gate_optimized   => G_use_gate_optimized,
          G_use_cascading        => G_use_cascading
        )
        port map (
          input  => f_input,
          output => f_output
        );

      -- AND Gate array
      -- generates each bit of the decoder result
      -- see block diagram
      coarse : for i in (c - 1) downto 0 generate -- generate columns

        fine : for j in (f - 1) downto 0 generate -- generate rows
          output((f * i) + j) <= c_output(i) and f_output(j);
        end generate fine;

      end generate coarse;

    else generate -- [G_use_cascading] is true

      -- cascaded decoders are generated recursively from the outside (final level) in

      -- * Configuration "Variables"

      function calc_liw (i: natural) return natural is

        variable prod     : real;
        variable exponent : real;

      begin

        prod := real(G_n);

        if (i > 1) then

          for j in 1 to (i - 1) loop

            prod := prod * (real(1) / calc_liw(j));

          end loop;

        end if;

        exponent := round(prod ** (real(1) / real(G_max_lvls - i + 1)));

        return natural(round(2 ** ceil(log2(exponent))));

      end function;

      constant liw_max : natural := calc_liw(G_max_lvls); -- L_m

      constant rem_in_width : natural := G_n / liw_max;

      -- output for the gestalt sub-decoder consisting of the remaining levels: 1 through [G_max_lvls] - 1
      signal rem_input  : std_logic_vector(lg(rem_in_width) - 1 downto 0);
      signal rem_output : std_logic_vector(rem_in_width - 1 downto 0);

      -- input for the final sub-decoder in the cascade
      signal l_max_input  : std_logic_vector(lg(liw_max) - 1 downto 0);
      signal l_max_output : std_logic_vector(liw_max - 1 downto 0);

    begin

      rem_input   <= input(G_lg_n - 1 downto lg(liw_max));
      l_max_input <= input(lg(liw_max) - 1 downto 0);

      dc_rem : ml_decoder
        generic map (
          G_n                    => rem_in_width,
          G_lg_n                 => lg(rem_in_width),
          G_max_lvls             => (G_max_lvls - 1),
          G_use_gate_optimized   => G_use_gate_optimized,
          G_use_cascading        => true
        )
        port map (
          input  => rem_input,
          output => rem_output
        );

      dc_l_max : ml_decoder
        generic map (
          G_n                    => liw_max,
          G_lg_n                 => lg(liw_max),
          G_max_lvls             => 1,
          G_use_gate_optimized   => G_use_gate_optimized,
          G_use_cascading        => false
        )
        port map (
          input  => l_max_input,
          output => l_max_output
        );

      -- AND Gate array
      -- generates each bit of the decoder result
      -- see block diagram
      arr_rem : for i in (rem_in_width - 1) downto 0 generate

        arr_l_max : for j in (liw_max - 1) downto 0 generate
          output((liw_max * i) + j) <= rem_output(i) and l_max_output(j);
        end generate arr_l_max;

      end generate arr_rem;

    end generate determine_encoder_type;

  else generate -- generate base level

    use_gate_optimized :
    if G_use_gate_optimized and (G_n = 4 or G_n = 8 or G_n = 16 or G_n = 32) generate
      -- This condition explicitly declares input widths in the case of inputs that are
      -- not powers of 2 causing synthesis to fail where the function-based option may "succeed".

      -- * Configuration "Variables"
      constant f    : natural := natural(round(2 ** ceil(log2(sqrt(real(G_n))))));  -- fine decoder output width
      constant lg_f : natural := lg(f);                                             -- fine decoder input width
      constant c    : natural := G_n / f;                                           -- coarse decoder output width
      constant lg_c : natural := lg(c);                                             -- coarse decoder input width

      signal c_input  : std_logic_vector(lg_c - 1 downto 0);  -- coarse decoder input
      signal c_output : std_logic_vector(c - 1 downto 0);     -- coarse decoder output
      signal f_input  : std_logic_vector(lg_f - 1 downto 0);  -- fine decoder input
      signal f_output : std_logic_vector(f - 1 downto 0);     -- fine decoder output      

    begin

      -- note that gate-level decoder boolean expressions correspond 
      --  to binary representation of a particular input value

      gate_lvl_dec :
      if (G_n = 32) generate -- 5:32 decoder
        
        c_output(3) <= input(4) and input(3);
        c_output(2) <= input(4) and not input(3);
        c_output(1) <= not input(4) and input(3);
        c_output(0) <= not input(4) and not input(3);

        f_output(7) <= input(2) and input(1) and input(0);
        f_output(6) <= input(2) and input(1) and not input(0);
        f_output(5) <= input(2) and not input(1) and input(0);
        f_output(4) <= input(2) and not input(1) and not input(0);
        f_output(3) <= not input(2) and input(1) and input(0);
        f_output(2) <= not input(2) and input(1) and not input(0);
        f_output(1) <= not input(2) and not input(1) and input(0);
        f_output(0) <= not input(2) and not input(1) and not input(0);
         
      elsif (G_n = 16) generate -- 4:16 decoder

        c_output(3) <= input(3) and input(2);
        c_output(2) <= input(3) and not input(2);
        c_output(1) <= not input(3) and input(2);
        c_output(0) <= not input(3) and not input(2);

        f_output(3) <= input(1) and input(0);
        f_output(2) <= input(1) and not input(0);
        f_output(1) <= not input(1) and input(0);
        f_output(0) <= not input(1) and not input(0);

      elsif (G_n = 8) generate -- 3:8 decoder

        c_output(1) <= input(2);
        c_output(0) <= not input(2);

        f_output(3) <= input(1) and input(0);
        f_output(2) <= input(1) and not input(0);
        f_output(1) <= not input(1) and input(0);
        f_output(0) <= not input(1) and not input(0);

      else generate -- 2:4 decoder

        c_output(1) <= input(1);
        c_output(0) <= not input(1);

        f_output(1) <= input(0);
        f_output(0) <= not input(0);

      end generate gate_lvl_dec;

      -- AND Gate array
      -- generates each bit of the decoder result
      -- see block diagram
      gld_coarse : for i in (c - 1) downto 0 generate -- generate columns

        gld_fine : for j in (f - 1) downto 0 generate -- generate rows
          output((f * i) + j) <= c_output(i) and f_output(j);
        end generate gld_fine;

      end generate gld_coarse;

    else generate -- generate function-based single-level decoder

      decoder : process (input) begin
        output <= (others => '0');

        output(natural(to_integer(unsigned(input)))) <= '1';
      end process;

    end generate use_gate_optimized;

  end generate determine_level;

end architecture behavioral;
