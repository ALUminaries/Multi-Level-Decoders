library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity decoder_262144 is
generic(
  g_n:      integer := 262144;  -- Input (multiplier) length is n
  g_log2n:  integer := 18;  -- Base 2 Logarithm of input length n; i.e., output length
  g_q:      integer := 512;  -- q is the least power of 2 greater than sqrt(n); i.e., 2^(ceil(log_2(sqrt(n)))
  g_log2q:  integer := 9;  -- Base 2 Logarithm of q
  g_k:      integer := 512;  -- k is defined as n/q, if n is a perfect square, then k = sqrt(n) = q
  g_log2k:  integer := 9  -- Base 2 Logarithm of k
);
port(
  input: in std_logic_vector(g_log2n - 1 downto 0); -- value to decode, i.e., shift amount for multiplication)
  output: out std_logic_vector(g_n - 1 downto 0) -- decoded result (C_i)
);
end decoder_262144;

architecture behavioral of decoder_262144 is

signal col: std_logic_vector(g_k - 1 downto 0); -- column/coarse decoder, handles log2k most significant bits of input
signal row: std_logic_vector(g_q - 1 downto 0); -- row/fine decoder, handles log2q least significant bits of input
signal result: std_logic_vector(g_n - 1 downto 0); -- result of decoding, i.e., 2^{input}

begin
-- Decoding corresponds to binary representation of given portions of shift

col(511) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(510) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(509) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(508) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(507) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(506) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(505) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(504) <= input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(503) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(502) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(501) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(500) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(499) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(498) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(497) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(496) <= input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(495) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(494) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(493) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(492) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(491) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(490) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(489) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(488) <= input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(487) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(486) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(485) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(484) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(483) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(482) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(481) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(480) <= input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(479) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(478) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(477) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(476) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(475) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(474) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(473) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(472) <= input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(471) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(470) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(469) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(468) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(467) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(466) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(465) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(464) <= input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(463) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(462) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(461) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(460) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(459) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(458) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(457) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(456) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(455) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(454) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(453) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(452) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(451) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(450) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(449) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(448) <= input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(447) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(446) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(445) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(444) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(443) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(442) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(441) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(440) <= input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(439) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(438) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(437) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(436) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(435) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(434) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(433) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(432) <= input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(431) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(430) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(429) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(428) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(427) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(426) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(425) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(424) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(423) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(422) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(421) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(420) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(419) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(418) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(417) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(416) <= input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(415) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(414) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(413) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(412) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(411) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(410) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(409) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(408) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(407) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(406) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(405) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(404) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(403) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(402) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(401) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(400) <= input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(399) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(398) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(397) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(396) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(395) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(394) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(393) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(392) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(391) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(390) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(389) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(388) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(387) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(386) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(385) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(384) <= input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(383) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(382) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(381) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(380) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(379) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(378) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(377) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(376) <= input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(375) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(374) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(373) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(372) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(371) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(370) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(369) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(368) <= input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(367) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(366) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(365) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(364) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(363) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(362) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(361) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(360) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(359) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(358) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(357) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(356) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(355) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(354) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(353) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(352) <= input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(351) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(350) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(349) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(348) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(347) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(346) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(345) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(344) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(343) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(342) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(341) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(340) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(339) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(338) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(337) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(336) <= input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(335) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(334) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(333) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(332) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(331) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(330) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(329) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(328) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(327) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(326) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(325) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(324) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(323) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(322) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(321) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(320) <= input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(319) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(318) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(317) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(316) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(315) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(314) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(313) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(312) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(311) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(310) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(309) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(308) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(307) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(306) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(305) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(304) <= input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(303) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(302) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(301) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(300) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(299) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(298) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(297) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(296) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(295) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(294) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(293) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(292) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(291) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(290) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(289) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(288) <= input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(287) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(286) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(285) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(284) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(283) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(282) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(281) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(280) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(279) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(278) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(277) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(276) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(275) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(274) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(273) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(272) <= input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(271) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(270) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(269) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(268) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(267) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(266) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(265) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(264) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(263) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(262) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(261) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(260) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(259) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(258) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(257) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(256) <= input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(255) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(254) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(253) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(252) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(251) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(250) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(249) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(248) <= not input(17) and input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(247) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(246) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(245) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(244) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(243) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(242) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(241) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(240) <= not input(17) and input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(239) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(238) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(237) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(236) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(235) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(234) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(233) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(232) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(231) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(230) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(229) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(228) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(227) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(226) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(225) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(224) <= not input(17) and input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(223) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(222) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(221) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(220) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(219) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(218) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(217) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(216) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(215) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(214) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(213) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(212) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(211) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(210) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(209) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(208) <= not input(17) and input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(207) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(206) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(205) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(204) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(203) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(202) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(201) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(200) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(199) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(198) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(197) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(196) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(195) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(194) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(193) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(192) <= not input(17) and input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(191) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(190) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(189) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(188) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(187) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(186) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(185) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(184) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(183) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(182) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(181) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(180) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(179) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(178) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(177) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(176) <= not input(17) and input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(175) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(174) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(173) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(172) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(171) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(170) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(169) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(168) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(167) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(166) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(165) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(164) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(163) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(162) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(161) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(160) <= not input(17) and input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(159) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(158) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(157) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(156) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(155) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(154) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(153) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(152) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(151) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(150) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(149) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(148) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(147) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(146) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(145) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(144) <= not input(17) and input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(143) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(142) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(141) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(140) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(139) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(138) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(137) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(136) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(135) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(134) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(133) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(132) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(131) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(130) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(129) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(128) <= not input(17) and input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(127) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(126) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(125) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(124) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(123) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(122) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(121) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(120) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(119) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(118) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(117) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(116) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(115) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(114) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(113) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(112) <= not input(17) and not input(16) and input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(111) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(110) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(109) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(108) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(107) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(106) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(105) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(104) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(103) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(102) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(101) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(100) <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(99)  <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(98)  <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(97)  <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(96)  <= not input(17) and not input(16) and input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(95)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(94)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(93)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(92)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(91)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(90)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(89)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(88)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(87)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(86)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(85)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(84)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(83)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(82)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(81)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(80)  <= not input(17) and not input(16) and input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(79)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(78)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(77)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(76)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(75)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(74)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(73)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(72)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(71)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(70)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(69)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(68)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(67)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(66)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(65)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(64)  <= not input(17) and not input(16) and input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(63)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(62)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(61)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(60)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(59)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(58)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(57)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(56)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(55)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(54)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(53)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(52)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(51)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(50)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(49)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(48)  <= not input(17) and not input(16) and not input(15) and input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(47)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(46)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(45)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(44)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(43)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(42)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(41)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(40)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(39)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(38)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(37)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(36)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(35)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(34)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(33)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(32)  <= not input(17) and not input(16) and not input(15) and input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(31)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and input(9);
col(30)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9);
col(29)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9);
col(28)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9);
col(27)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9);
col(26)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9);
col(25)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9);
col(24)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(23)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9);
col(22)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9);
col(21)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9);
col(20)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(19)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9);
col(18)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(17)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(16)  <= not input(17) and not input(16) and not input(15) and not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9);
col(15)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9);
col(14)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9);
col(13)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9);
col(12)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9);
col(11)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9);
col(10)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9);
col(9)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9);
col(8)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9);
col(7)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9);
col(6)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9);
col(5)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9);
col(4)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9);
col(3)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9);
col(2)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9);
col(1)   <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9);
col(0)  <= not input(17) and not input(16) and not input(15) and not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9);

row(511) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(510) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(509) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(508) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(507) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(506) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(505) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(504) <= input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(503) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(502) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(501) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(500) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(499) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(498) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(497) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(496) <= input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(495) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(494) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(493) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(492) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(491) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(490) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(489) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(488) <= input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(487) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(486) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(485) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(484) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(483) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(482) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(481) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(480) <= input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(479) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(478) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(477) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(476) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(475) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(474) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(473) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(472) <= input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(471) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(470) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(469) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(468) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(467) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(466) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(465) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(464) <= input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(463) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(462) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(461) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(460) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(459) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(458) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(457) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(456) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(455) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(454) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(453) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(452) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(451) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(450) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(449) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(448) <= input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(447) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(446) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(445) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(444) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(443) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(442) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(441) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(440) <= input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(439) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(438) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(437) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(436) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(435) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(434) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(433) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(432) <= input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(431) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(430) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(429) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(428) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(427) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(426) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(425) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(424) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(423) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(422) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(421) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(420) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(419) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(418) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(417) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(416) <= input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(415) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(414) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(413) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(412) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(411) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(410) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(409) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(408) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(407) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(406) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(405) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(404) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(403) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(402) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(401) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(400) <= input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(399) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(398) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(397) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(396) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(395) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(394) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(393) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(392) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(391) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(390) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(389) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(388) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(387) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(386) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(385) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(384) <= input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(383) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(382) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(381) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(380) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(379) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(378) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(377) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(376) <= input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(375) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(374) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(373) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(372) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(371) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(370) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(369) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(368) <= input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(367) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(366) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(365) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(364) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(363) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(362) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(361) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(360) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(359) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(358) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(357) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(356) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(355) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(354) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(353) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(352) <= input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(351) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(350) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(349) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(348) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(347) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(346) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(345) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(344) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(343) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(342) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(341) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(340) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(339) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(338) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(337) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(336) <= input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(335) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(334) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(333) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(332) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(331) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(330) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(329) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(328) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(327) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(326) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(325) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(324) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(323) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(322) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(321) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(320) <= input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(319) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(318) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(317) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(316) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(315) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(314) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(313) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(312) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(311) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(310) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(309) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(308) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(307) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(306) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(305) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(304) <= input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(303) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(302) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(301) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(300) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(299) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(298) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(297) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(296) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(295) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(294) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(293) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(292) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(291) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(290) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(289) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(288) <= input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(287) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(286) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(285) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(284) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(283) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(282) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(281) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(280) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(279) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(278) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(277) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(276) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(275) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(274) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(273) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(272) <= input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(271) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(270) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(269) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(268) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(267) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(266) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(265) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(264) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(263) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(262) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(261) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(260) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(259) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(258) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(257) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(256) <= input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(255) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(254) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(253) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(252) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(251) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(250) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(249) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(248) <= not input(8) and input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(247) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(246) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(245) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(244) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(243) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(242) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(241) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(240) <= not input(8) and input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(239) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(238) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(237) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(236) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(235) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(234) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(233) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(232) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(231) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(230) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(229) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(228) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(227) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(226) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(225) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(224) <= not input(8) and input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(223) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(222) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(221) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(220) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(219) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(218) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(217) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(216) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(215) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(214) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(213) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(212) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(211) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(210) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(209) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(208) <= not input(8) and input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(207) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(206) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(205) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(204) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(203) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(202) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(201) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(200) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(199) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(198) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(197) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(196) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(195) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(194) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(193) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(192) <= not input(8) and input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(191) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(190) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(189) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(188) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(187) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(186) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(185) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(184) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(183) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(182) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(181) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(180) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(179) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(178) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(177) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(176) <= not input(8) and input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(175) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(174) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(173) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(172) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(171) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(170) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(169) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(168) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(167) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(166) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(165) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(164) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(163) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(162) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(161) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(160) <= not input(8) and input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(159) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(158) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(157) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(156) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(155) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(154) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(153) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(152) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(151) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(150) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(149) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(148) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(147) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(146) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(145) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(144) <= not input(8) and input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(143) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(142) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(141) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(140) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(139) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(138) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(137) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(136) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(135) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(134) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(133) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(132) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(131) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(130) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(129) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(128) <= not input(8) and input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(127) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(126) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(125) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(124) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(123) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(122) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(121) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(120) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(119) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(118) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(117) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(116) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(115) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(114) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(113) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(112) <= not input(8) and not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(111) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(110) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(109) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(108) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(107) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(106) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(105) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(104) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(103) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(102) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(101) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(100) <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(99)  <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(98)  <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(97)  <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(96)  <= not input(8) and not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(95)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(94)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(93)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(92)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(91)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(90)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(89)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(88)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(87)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(86)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(85)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(84)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(83)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(82)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(81)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(80)  <= not input(8) and not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(79)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(78)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(77)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(76)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(75)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(74)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(73)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(72)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(71)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(70)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(69)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(68)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(67)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(66)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(65)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(64)  <= not input(8) and not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(63)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(62)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(61)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(60)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(59)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(58)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(57)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(56)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(55)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(54)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(53)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(52)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(51)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(50)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(49)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(48)  <= not input(8) and not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(47)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(46)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(45)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(44)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(43)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(42)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(41)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(40)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(39)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(38)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(37)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(36)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(35)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(34)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(33)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(32)  <= not input(8) and not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(31)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(30)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(29)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(28)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(27)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(26)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(25)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(24)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(23)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(22)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(21)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(20)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(19)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(18)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(17)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(16)  <= not input(8) and not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(15)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(14)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(13)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(12)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(11)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(10)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(9)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(8)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(7)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(6)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(5)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(4)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(3)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(2)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(1)   <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(0)  <= not input(8) and not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);


-- generates each bit of the decoder result
-- see two-level decoder block diagram
coarse: for i in g_k - 1 downto 0 generate -- generate columns
  fine: for j in g_q - 1 downto 0 generate -- generate rows
    result((g_q * i) + j) <= col(i) and row(j);
  end generate fine;
end generate coarse;

output <= result;
end;