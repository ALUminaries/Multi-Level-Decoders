library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity decoder_32768 is
generic(
  g_n:      integer := 32768;  -- Input (multiplier) length is n
  g_log2n:  integer := 15;  -- Base 2 Logarithm of input length n; i.e., output length
  g_q:      integer := 256;  -- q is the least power of 2 greater than sqrt(n); i.e., 2^(ceil(log_2(sqrt(n)))
  g_log2q:  integer := 8;  -- Base 2 Logarithm of q
  g_k:      integer := 128;  -- k is defined as n/q, if n is a perfect square, then k = sqrt(n) = q
  g_log2k:  integer := 7  -- Base 2 Logarithm of k
);
port(
  input: in std_logic_vector(g_log2n - 1 downto 0); -- value to decode, i.e., shift amount for multiplication)
  output: out std_logic_vector(g_n - 1 downto 0) -- decoded result (C_i)
);
end decoder_32768;

architecture behavioral of decoder_32768 is

signal col: std_logic_vector(g_k - 1 downto 0); -- column/coarse decoder, handles log2k most significant bits of input
signal row: std_logic_vector(g_q - 1 downto 0); -- row/fine decoder, handles log2q least significant bits of input
signal result: std_logic_vector(g_n - 1 downto 0); -- result of decoding, i.e., 2^{input}

begin
-- Decoding corresponds to binary representation of given portions of shift

col(127) <= input(14) and input(13) and input(12) and input(11) and input(10) and input(9) and input(8);
col(126) <= input(14) and input(13) and input(12) and input(11) and input(10) and input(9) and not input(8);
col(125) <= input(14) and input(13) and input(12) and input(11) and input(10) and not input(9) and input(8);
col(124) <= input(14) and input(13) and input(12) and input(11) and input(10) and not input(9) and not input(8);
col(123) <= input(14) and input(13) and input(12) and input(11) and not input(10) and input(9) and input(8);
col(122) <= input(14) and input(13) and input(12) and input(11) and not input(10) and input(9) and not input(8);
col(121) <= input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9) and input(8);
col(120) <= input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(119) <= input(14) and input(13) and input(12) and not input(11) and input(10) and input(9) and input(8);
col(118) <= input(14) and input(13) and input(12) and not input(11) and input(10) and input(9) and not input(8);
col(117) <= input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9) and input(8);
col(116) <= input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(115) <= input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9) and input(8);
col(114) <= input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(113) <= input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(112) <= input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(111) <= input(14) and input(13) and not input(12) and input(11) and input(10) and input(9) and input(8);
col(110) <= input(14) and input(13) and not input(12) and input(11) and input(10) and input(9) and not input(8);
col(109) <= input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9) and input(8);
col(108) <= input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9) and not input(8);
col(107) <= input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9) and input(8);
col(106) <= input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9) and not input(8);
col(105) <= input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9) and input(8);
col(104) <= input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(103) <= input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9) and input(8);
col(102) <= input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9) and not input(8);
col(101) <= input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9) and input(8);
col(100) <= input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(99)  <= input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9) and input(8);
col(98)  <= input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(97)  <= input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(96)  <= input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(95)  <= input(14) and not input(13) and input(12) and input(11) and input(10) and input(9) and input(8);
col(94)  <= input(14) and not input(13) and input(12) and input(11) and input(10) and input(9) and not input(8);
col(93)  <= input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9) and input(8);
col(92)  <= input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9) and not input(8);
col(91)  <= input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9) and input(8);
col(90)  <= input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9) and not input(8);
col(89)  <= input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9) and input(8);
col(88)  <= input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(87)  <= input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9) and input(8);
col(86)  <= input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9) and not input(8);
col(85)  <= input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9) and input(8);
col(84)  <= input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(83)  <= input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9) and input(8);
col(82)  <= input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(81)  <= input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(80)  <= input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(79)  <= input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9) and input(8);
col(78)  <= input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9) and not input(8);
col(77)  <= input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9) and input(8);
col(76)  <= input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9) and not input(8);
col(75)  <= input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9) and input(8);
col(74)  <= input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9) and not input(8);
col(73)  <= input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9) and input(8);
col(72)  <= input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(71)  <= input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9) and input(8);
col(70)  <= input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9) and not input(8);
col(69)  <= input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9) and input(8);
col(68)  <= input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(67)  <= input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9) and input(8);
col(66)  <= input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(65)  <= input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(64)  <= input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(63)  <= not input(14) and input(13) and input(12) and input(11) and input(10) and input(9) and input(8);
col(62)  <= not input(14) and input(13) and input(12) and input(11) and input(10) and input(9) and not input(8);
col(61)  <= not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9) and input(8);
col(60)  <= not input(14) and input(13) and input(12) and input(11) and input(10) and not input(9) and not input(8);
col(59)  <= not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9) and input(8);
col(58)  <= not input(14) and input(13) and input(12) and input(11) and not input(10) and input(9) and not input(8);
col(57)  <= not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9) and input(8);
col(56)  <= not input(14) and input(13) and input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(55)  <= not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9) and input(8);
col(54)  <= not input(14) and input(13) and input(12) and not input(11) and input(10) and input(9) and not input(8);
col(53)  <= not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9) and input(8);
col(52)  <= not input(14) and input(13) and input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(51)  <= not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9) and input(8);
col(50)  <= not input(14) and input(13) and input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(49)  <= not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(48)  <= not input(14) and input(13) and input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(47)  <= not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9) and input(8);
col(46)  <= not input(14) and input(13) and not input(12) and input(11) and input(10) and input(9) and not input(8);
col(45)  <= not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9) and input(8);
col(44)  <= not input(14) and input(13) and not input(12) and input(11) and input(10) and not input(9) and not input(8);
col(43)  <= not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9) and input(8);
col(42)  <= not input(14) and input(13) and not input(12) and input(11) and not input(10) and input(9) and not input(8);
col(41)  <= not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9) and input(8);
col(40)  <= not input(14) and input(13) and not input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(39)  <= not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9) and input(8);
col(38)  <= not input(14) and input(13) and not input(12) and not input(11) and input(10) and input(9) and not input(8);
col(37)  <= not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9) and input(8);
col(36)  <= not input(14) and input(13) and not input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(35)  <= not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9) and input(8);
col(34)  <= not input(14) and input(13) and not input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(33)  <= not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(32)  <= not input(14) and input(13) and not input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(31)  <= not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9) and input(8);
col(30)  <= not input(14) and not input(13) and input(12) and input(11) and input(10) and input(9) and not input(8);
col(29)  <= not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9) and input(8);
col(28)  <= not input(14) and not input(13) and input(12) and input(11) and input(10) and not input(9) and not input(8);
col(27)  <= not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9) and input(8);
col(26)  <= not input(14) and not input(13) and input(12) and input(11) and not input(10) and input(9) and not input(8);
col(25)  <= not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9) and input(8);
col(24)  <= not input(14) and not input(13) and input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(23)  <= not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9) and input(8);
col(22)  <= not input(14) and not input(13) and input(12) and not input(11) and input(10) and input(9) and not input(8);
col(21)  <= not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9) and input(8);
col(20)  <= not input(14) and not input(13) and input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(19)  <= not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9) and input(8);
col(18)  <= not input(14) and not input(13) and input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(17)  <= not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(16)  <= not input(14) and not input(13) and input(12) and not input(11) and not input(10) and not input(9) and not input(8);
col(15)  <= not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9) and input(8);
col(14)  <= not input(14) and not input(13) and not input(12) and input(11) and input(10) and input(9) and not input(8);
col(13)  <= not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9) and input(8);
col(12)  <= not input(14) and not input(13) and not input(12) and input(11) and input(10) and not input(9) and not input(8);
col(11)  <= not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9) and input(8);
col(10)  <= not input(14) and not input(13) and not input(12) and input(11) and not input(10) and input(9) and not input(8);
col(9)   <= not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9) and input(8);
col(8)   <= not input(14) and not input(13) and not input(12) and input(11) and not input(10) and not input(9) and not input(8);
col(7)   <= not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9) and input(8);
col(6)   <= not input(14) and not input(13) and not input(12) and not input(11) and input(10) and input(9) and not input(8);
col(5)   <= not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9) and input(8);
col(4)   <= not input(14) and not input(13) and not input(12) and not input(11) and input(10) and not input(9) and not input(8);
col(3)   <= not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9) and input(8);
col(2)   <= not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and input(9) and not input(8);
col(1)   <= not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9) and input(8);
col(0)  <= not input(14) and not input(13) and not input(12) and not input(11) and not input(10) and not input(9) and not input(8);

row(255) <= input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(254) <= input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(253) <= input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(252) <= input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(251) <= input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(250) <= input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(249) <= input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(248) <= input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(247) <= input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(246) <= input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(245) <= input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(244) <= input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(243) <= input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(242) <= input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(241) <= input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(240) <= input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(239) <= input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(238) <= input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(237) <= input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(236) <= input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(235) <= input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(234) <= input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(233) <= input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(232) <= input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(231) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(230) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(229) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(228) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(227) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(226) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(225) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(224) <= input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(223) <= input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(222) <= input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(221) <= input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(220) <= input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(219) <= input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(218) <= input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(217) <= input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(216) <= input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(215) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(214) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(213) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(212) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(211) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(210) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(209) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(208) <= input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(207) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(206) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(205) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(204) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(203) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(202) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(201) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(200) <= input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(199) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(198) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(197) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(196) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(195) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(194) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(193) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(192) <= input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(191) <= input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(190) <= input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(189) <= input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(188) <= input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(187) <= input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(186) <= input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(185) <= input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(184) <= input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(183) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(182) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(181) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(180) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(179) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(178) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(177) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(176) <= input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(175) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(174) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(173) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(172) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(171) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(170) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(169) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(168) <= input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(167) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(166) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(165) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(164) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(163) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(162) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(161) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(160) <= input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(159) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(158) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(157) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(156) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(155) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(154) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(153) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(152) <= input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(151) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(150) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(149) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(148) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(147) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(146) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(145) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(144) <= input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(143) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(142) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(141) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(140) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(139) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(138) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(137) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(136) <= input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(135) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(134) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(133) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(132) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(131) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(130) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(129) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(128) <= input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(127) <= not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(126) <= not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(125) <= not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(124) <= not input(7) and input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(123) <= not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(122) <= not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(121) <= not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(120) <= not input(7) and input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(119) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(118) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(117) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(116) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(115) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(114) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(113) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(112) <= not input(7) and input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(111) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(110) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(109) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(108) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(107) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(106) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(105) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(104) <= not input(7) and input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(103) <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(102) <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(101) <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(100) <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(99)  <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(98)  <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(97)  <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(96)  <= not input(7) and input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(95)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(94)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(93)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(92)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(91)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(90)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(89)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(88)  <= not input(7) and input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(87)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(86)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(85)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(84)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(83)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(82)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(81)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(80)  <= not input(7) and input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(79)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(78)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(77)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(76)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(75)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(74)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(73)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(72)  <= not input(7) and input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(71)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(70)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(69)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(68)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(67)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(66)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(65)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(64)  <= not input(7) and input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(63)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(62)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(61)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(60)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(59)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(58)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(57)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(56)  <= not input(7) and not input(6) and input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(55)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(54)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(53)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(52)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(51)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(50)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(49)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(48)  <= not input(7) and not input(6) and input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(47)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(46)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(45)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(44)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(43)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(42)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(41)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(40)  <= not input(7) and not input(6) and input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(39)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(38)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(37)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(36)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(35)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(34)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(33)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(32)  <= not input(7) and not input(6) and input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(31)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and input(0);
row(30)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and input(1) and not input(0);
row(29)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and input(0);
row(28)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and input(2) and not input(1) and not input(0);
row(27)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and input(0);
row(26)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and input(1) and not input(0);
row(25)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and input(0);
row(24)  <= not input(7) and not input(6) and not input(5) and input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(23)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and input(0);
row(22)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and input(1) and not input(0);
row(21)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and input(0);
row(20)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(19)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and input(0);
row(18)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(17)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(16)  <= not input(7) and not input(6) and not input(5) and input(4) and not input(3) and not input(2) and not input(1) and not input(0);
row(15)  <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and input(0);
row(14)  <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and input(1) and not input(0);
row(13)  <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and input(0);
row(12)  <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and input(2) and not input(1) and not input(0);
row(11)  <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and input(0);
row(10)  <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and input(1) and not input(0);
row(9)   <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and input(0);
row(8)   <= not input(7) and not input(6) and not input(5) and not input(4) and input(3) and not input(2) and not input(1) and not input(0);
row(7)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and input(0);
row(6)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and input(1) and not input(0);
row(5)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and input(0);
row(4)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and input(2) and not input(1) and not input(0);
row(3)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and input(0);
row(2)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and input(1) and not input(0);
row(1)   <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and input(0);
row(0)  <= not input(7) and not input(6) and not input(5) and not input(4) and not input(3) and not input(2) and not input(1) and not input(0);


-- generates each bit of the decoder result
-- see two-level decoder block diagram
coarse: for i in g_k - 1 downto 0 generate -- generate columns
  fine: for j in g_q - 1 downto 0 generate -- generate rows
    result((g_q * i) + j) <= col(i) and row(j);
  end generate fine;
end generate coarse;

output <= result;
end;